package merger;
import FixedPoint::*;
import FIFO::*;
import FIFOF::*;
import datatypes::*;
import SpecialFIFOs:: * ;
import Real::*;
import Vector::*;

#define REPL 128


#define BWIDTH0 8
#define BWIDTH1 16
#define BWIDTH2 24
#define BWIDTH7 24


interface Merge;
        method Action put(Vector#(REPL, DataType) datas);
        method ActionValue#(Vector#(REPL, Vector#(3,Bit#(BWIDTH7)))) get;
	method Action configure(UInt#(4) a, Bit#(8) m, UInt#(6) wx);	
endinterface

(*synthesize*)
module mkMerge(Merge);
Reg#(UInt#(4))  kernel   <- mkReg(0);
Reg#(Bit#(8))   mx       <- mkReg(0);
Reg#(UInt#(6)) cx        <- mkReg(0);
Reg#(UInt#(6)) width     <- mkReg(16);

Reg#(Bit#(BWIDTH0))  _L1[REPL];
Reg#(Bit#(BWIDTH1))  _L2[REPL];
Reg#(Bit#(BWIDTH2))  _L3[REPL];
Reg#(Bit#(BWIDTH2))  _L9[3*REPL];


for(int i=0;i<REPL;i=i+1) begin
	_L1[i]   <- mkReg(0);
	_L2[i]   <- mkReg(0);
	_L3[i]   <- mkReg(0);
end

for(int i=0;i<3*REPL;i=i+1) 
	_L9[i]   <- mkReg(0);


FIFOF#(Bit#(1)) p0 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p1 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p2 <- mkPipelineFIFOF;
FIFOF#(Bit#(1)) p3 <- mkPipelineFIFOF;

	//###########################################################


	for(int i=0;i< REPL-1; i = i + 1) begin 
	rule _Q1;
		Bit#(BWIDTH1) x1    = extend(_L1[i]);
		Bit#(BWIDTH1) x2    = extend(_L1[i+1]);
		Bit#(BWIDTH1) y     = (x1 << 8) | x2;
		_L2[i] <= y;	
	endrule

	
	rule _Q2;
		Bit#(BWIDTH2) x1    = extend(_L2[i]);
		Bit#(BWIDTH2) x2    = extend(_L2[i+1]);
		Bit#(BWIDTH2) y     = (x1 << 8) | x2;
		_L3[i] <= y;	
        endrule
	end	
	//################################################
	
    	rule _activate1;
		p0.deq;
		p1.enq(1);
    	endrule

   	rule _activate2;
		p1.deq;
		p2.enq(1);
    	endrule
	//################################################
	

	rule coalesce;
		p2.deq;
		for(int i=0;i<REPL; i = i + 1) begin
			Vector#(3,DataType) mx = unpack(_L3[i]);
			for(int j=0;j<3;j=j+1)
                	_L9[i*3+j]          <= (_L9[i*3+j] << 8) | zeroExtend(pack(mx[j]));
		end
		if (cx >= zeroExtend(kernel-1))
			p3.enq(1);

		if (cx == width-1)
                        cx <= 0;
                else
                        cx <= cx + 1;
	endrule
		
        method Action put(Vector#(REPL, DataType) datas);
		for(int i = 0; i <REPL; i = i + 1)
			_L1[i] <= pack(datas[i]);	
		p0.enq(1);
	endmethod
	
        method ActionValue#(Vector#(REPL, Vector#(3,Bit#(BWIDTH7)))) get;
		p3.deq;
		Vector#(REPL, Vector#(3,Bit#(BWIDTH7))) out = newVector;
		for(int i=0;i<REPL; i = i + 1)
			for(int j=0;j<3;j=j+1)
			out[i][j] = _L9[i*3+j];
		return out;
	endmethod
	
	method Action configure(UInt#(4) a, Bit#(8) m, UInt#(6) wx);	
			kernel  <= 3;
			mx 	<= m;
			width   <= wx;
	endmethod
	
endmodule
endpackage
